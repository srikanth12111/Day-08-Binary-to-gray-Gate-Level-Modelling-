`timescale 1ns / 1ps
module binary_to_gray_tb;
reg b1,b2,b3,b4;
wire g1,g2,g3,g4;
binary_to_gray DUT(.b1(b1),.b2(b2),.b3(b3),.b4(b4),.g1(g1),.g2(g2),.g3(g3),.g4(g4));
initial
begin
b1 = 0;b2 = 0;b3 = 0;b4 = 0;
#100
#100 b1 = 0; b2 = 0; b3 = 0; b4 = 1;
#100 b1 = 0; b2 = 0; b3 = 1; b4 = 0;
#100 b1 = 0; b2 = 0; b3 = 1; b4 = 1;
#100 b1 = 0; b2 = 1; b3 = 0; b4 = 0;
#100 b1 = 0; b2 = 1; b3 = 0; b4 = 1;
#100 b1 = 0; b2 = 1; b3 = 1; b4 = 0;
#100 b1 = 0; b2 = 1; b3 = 1; b4 = 1;
#100 b1 = 1; b2 = 0; b3 = 0; b4 = 0;
#100 b1 = 1; b2 = 0; b3 = 0; b4 = 1;
#100 b1 = 1; b2 = 0; b3 = 1; b4 = 0;
#100 b1 = 1; b2 = 0; b3 = 1; b4 = 1;
#100 b1 = 1; b2 = 1; b3 = 0; b4 = 0;
#100 b1 = 1; b2 = 1; b3 = 0; b4 = 1;
#100 b1 = 1; b2 = 1; b3 = 1; b4 = 0;
#100 b1 = 1; b2 = 1; b3 = 1; b4 = 1;
end
endmodule
